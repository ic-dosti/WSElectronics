** Profile: "SCHEMATIC1-FFT"  [ C:\Users\useroot\Documents\GitHub\DOSTI\ExperimentalProjects\Cadence Allegro\LT1167\lt1167_pspice-pspicefiles\schematic1\fft.sim ] 

** Creating circuit file "FFT.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\useroot\Documents\Cadence\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
